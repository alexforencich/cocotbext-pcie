
`resetall
`timescale 1 ns / 1 ps
`default_nettype none

module test_pcie;

endmodule

`resetall
